.title KiCad schematic
R12 OUT Net-_R12-Pad2_ 100k
XU1 OUT Net-_R12-Pad2_ Net-_R1-Pad2_ +15V Net-_R13-Pad2_ Net-_R2-Pad2_ Net-_R13-Pad1_ Net-_R14-Pad1_ Net-_R3-Pad2_ Net-_R14-Pad2_ -15V Net-_R10-Pad1_ Net-_R4-Pad2_ Net-_R15-Pad1_ LM324c
XU2 Net-_R16-Pad1_ Net-_R11-Pad1_ Net-_R5-Pad2_ +15V NC_01 NC_02 NC_03 NC_04 NC_05 NC_06 -15V NC_07 NC_08 NC_09 LM324c
R16 Net-_R16-Pad1_ Net-_R11-Pad1_ 100k
R15 Net-_R15-Pad1_ Net-_R10-Pad1_ 100k
R14 Net-_R14-Pad1_ Net-_R14-Pad2_ 100k
R13 Net-_R13-Pad1_ Net-_R13-Pad2_ 100k
R6 Net-_R5-Pad2_ -15V 150k
R5 Net-_R4-Pad2_ Net-_R5-Pad2_ 47k
R11 Net-_R11-Pad1_ CV 10k
R4 Net-_R3-Pad2_ Net-_R4-Pad2_ 47k
R3 Net-_R2-Pad2_ Net-_R3-Pad2_ 47k
R10 Net-_R10-Pad1_ CV 10k
R9 Net-_R14-Pad2_ CV 10k
R8 Net-_R13-Pad2_ CV 10k
R7 Net-_R12-Pad2_ CV 10k
R2 Net-_R1-Pad2_ Net-_R2-Pad2_ 47k
R1 +15V Net-_R1-Pad2_ 150k
.end
