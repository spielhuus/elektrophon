.title KiCad schematic
R1 Net-_C1-Pad1_ GND 470k
C1 Net-_C1-Pad1_ IN 10u
XRV1 Net-_Q2-Pad1_ Net-_C5-Pad1_ Net-_R9-Pad2_ voltage_divider
R3 Net-_C3-Pad2_ GND 1k
C3 GND Net-_C3-Pad2_ 10u
R5 Net-_C4-Pad2_ GND 1.5k
C4 GND Net-_C4-Pad2_ 10u
C7 Net-_C7-Pad1_ +15V 47n
R8 Net-_C7-Pad1_ +15V 100k
C5 Net-_C5-Pad1_ Net-_C2-Pad1_ 2.2n
R7 Net-_Q2-Pad1_ Net-_C6-Pad1_ 1.2Meg
C6 Net-_C6-Pad1_ Net-_C2-Pad1_ 47n
R6 Net-_C2-Pad1_ Net-_C1-Pad1_ 2.2Meg
R4 Net-_C7-Pad1_ Net-_Q2-Pad1_ 47k
R2 +15V Net-_C2-Pad1_ 22k
C2 Net-_C2-Pad1_ Net-_C1-Pad1_ 1n
Q1 Net-_C2-Pad1_ Net-_C1-Pad1_ Net-_C3-Pad2_ BC547B
Q2 Net-_Q2-Pad1_ Net-_C6-Pad1_ Net-_C4-Pad2_ BC547B
R9 OUT Net-_R9-Pad2_ 100k
R10 GND OUT 20k
.end
