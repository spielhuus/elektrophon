.title KiCad schematic
R5 Net-_C1-Pad2_ Net-_Q1-Pad1_ 10k
R4 -15V Net-_Q2-Pad3_ 22k
R3 Net-_Q1-Pad3_ +15V 22k
R1 Net-_Q1-Pad2_ NC_01 27k
R2 Net-_Q1-Pad2_ GND 68k
R8 Net-_C1-Pad1_ Net-_C1-Pad2_ 120k
C1 Net-_C1-Pad1_ Net-_C1-Pad2_ 27p
C4 NC_02 Net-_C1-Pad1_ 680n
Q2 Net-_Q1-Pad1_ Net-_Q1-Pad2_ Net-_Q2-Pad3_ BC549
Q1 Net-_Q1-Pad1_ Net-_Q1-Pad2_ Net-_Q1-Pad3_ BC559
U1 GND Net-_C1-Pad2_ Net-_C1-Pad1_ TL074
.end
