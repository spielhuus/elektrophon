.title KiCad schematic
XU4 Net-_C3-Pad2_ Net-_C3-Pad1_ +5V GND 4069UB
C1 Net-_C1-Pad1_ IN 1u
XU1 Net-_C1-Pad1_ Net-_R2-Pad1_ +5V GND 4069UB
R2 Net-_R2-Pad1_ Net-_C1-Pad1_ 100k
R1 Net-_C2-Pad1_ Net-_C1-Pad1_ 100k
R3 Net-_R3-Pad1_ Net-_R2-Pad1_ 100k
XU2 Net-_R3-Pad1_ Net-_R4-Pad1_ +5V GND 4069UB
R4 Net-_R4-Pad1_ Net-_R3-Pad1_ 100k
XRV2 NC_01 Net-_C2-Pad2_ Net-_R5-Pad1_ voltage_divider_2
R5 Net-_R5-Pad1_ Net-_R4-Pad1_ 1k
XU3 Net-_C2-Pad2_ Net-_C2-Pad1_ +5V GND 4069UB
C2 Net-_C2-Pad1_ Net-_C2-Pad2_ 0.01u
XRV3 NC_02 Net-_C3-Pad2_ Net-_R6-Pad1_ voltage_divider_3
R6 Net-_R6-Pad1_ Net-_C2-Pad1_ 1k
C3 Net-_C3-Pad1_ Net-_C3-Pad2_ 0.01u
XRV1 NC_03 Net-_R3-Pad1_ Net-_C3-Pad1_ voltage_divider_1
C4 OUT Net-_C3-Pad1_ 1u
R7 GND OUT 1k
.end
