.title KiCad schematic
C3 GND -15V 10u
C2 +15V GND 10u
J1 -15V -15V +15V +15V GND GND GND GND +5V +5V IDC Header
IC1 -15V +15V RC4136
C4 +15V GND 0.1u
C5 GND -15V 0.1u
C7 +15V GND 0.1u
C8 GND -15V 0.1u
H1 MountingHole
H2 MountingHole
H3 MountingHole
H4 MountingHole
U2 -15V +15V SSM2040
J2 +15V -15V GND NC_01 NC_02 NC_03 NC_04 Conn_01x07_Female
C11 GND -15V 0.1u
C10 +15V GND 0.1u
C17 GND -15V 0.1u
C16 +15V GND 0.1u
U4 NC_05 NC_06 GND +15V NC_07 NC_08 -15V NC_09 LM4250
U6 NC_10 NC_11 NC_12 -15V NC_13 NC_14 +15V NC_15 LM4250
U1 Net-_RV1-Pad1_ Net-_RV1-Pad1_ Net-_R6-Pad1_ NC_16 GND Net-_R10-Pad2_ Net-_R10-Pad1_ NC_17 TL072
U3 Net-_Q1-Pad1_ Net-_R11-Pad1_ GND NC_18 NC_19 NC_20 NC_21 NC_22 TL072
U5 NC_23 NC_24 NC_25 NC_26 NC_27 NC_28 NC_29 NC_30 TL072
J3 GND Net-_J3-PadT_ NC_31 FM_IN
R6 Net-_R6-Pad1_ Net-_J3-PadT_ 10k
RV1 Net-_RV1-Pad1_ Net-_R11-Pad2_ Net-_R10-Pad1_ 47k
R10 Net-_R10-Pad1_ Net-_R10-Pad2_ 100k
R5 Net-_R10-Pad2_ Net-_J3-PadT_ 100k
R3 GND Net-_J3-PadT_ 220k
R11 Net-_R11-Pad1_ Net-_R11-Pad2_ 120k
R15 Net-_Q1-Pad1_ Net-_R11-Pad1_ 3k
Q1 Net-_Q1-Pad1_ Net-_Q1-Pad1_ NC_32 2N3904
RV2 +15V Net-_R4-Pad2_ Net-_R1-Pad2_ 100k
R1 -15V Net-_R1-Pad2_ 47k
R4 Net-_R11-Pad1_ Net-_R4-Pad2_ 162k
J4 GND Net-_J4-PadT_ NC_33 CV_IN
J5 GND Net-_J5-PadT_ NC_34 INPUT
R7 Net-_R11-Pad1_ Net-_J4-PadT_ 100k
R14 Net-_R11-Pad1_ +15V 100k
R8 NC_35 Net-_J5-PadT_ 470k
R12 Net-_R12-Pad1_ NC_36 47k
R13 GND Net-_R12-Pad1_ 1k
R9 NC_37 NC_38 27k
RV3 NC_39 NC_40 Net-_R2-Pad2_ 100k
R2 GND Net-_R2-Pad2_ 100
.end
