.title KiCad schematic
Q9 Net-_Q10-Pad2_ Net-_Q9-Pad2_ Net-_C12-Pad1_ BC846B
Q10 Net-_C12-Pad1_ Net-_Q10-Pad2_ +15V BC556B
R26 Net-_Q9-Pad2_ Net-_C11-Pad1_ 10k
R25 Net-_C12-Pad2_ Net-_C11-Pad1_ 15k
C11 Net-_C11-Pad1_ GND 22n
C12 Net-_C12-Pad1_ Net-_C12-Pad2_ 220n
R24 Net-_C12-Pad2_ NC_01 15k
R27 GND Net-_C12-Pad1_ 1.5k
C13 OUT Net-_C12-Pad1_ 100u
R28 GND OUT 10k
.end
