.title KiCad schematic
.include ../../../lib/spice/cmos/CD4069UB-hex.lib
.include ../../../lib/spice/diode/1N4148.mod
.include 'UBE Screamer.cir'
.control
* Save only the output values
save v(OUT)
* 44100Hz sampling frequency
tran 22.675u 6
wrdata build/output v(OUT)
* you can use output.data as input for scripts
.endc
.subckt voltage_divider_1 n1 n2 n3
R1 n1 n2 499kOhm
R2 n2 n3 1kOhm
.ends voltage_divider_1

.subckt voltage_divider_2 n1 n2 n3
R1 n1 n2 1.0kOhm
R2 n2 n3 500.0kOhm
.ends voltage_divider_2
V1 +5V 0 DC 5
a1 %v([IN]) filesrc

.model filesrc filesource (file="build/input.spice" amploffset=[0] amplscale=[5]
+                          timeoffset=0 timescale=1
+                          timerelative=false amplstep=false)

.end
.measure tran ymax MAX v(OUT) from=0m to=30m
.measure tran ymax RMS v(OUT) from=0m to=30m

