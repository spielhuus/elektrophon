.title KiCad schematic
Q2 Net-_Q2-Pad1_ Net-_C6-Pad1_ Net-_C4-Pad2_ BC547B
Q1 Net-_C2-Pad1_ Net-_C1-Pad1_ Net-_C3-Pad2_ BC547B
R1 Net-_C1-Pad1_ GND 470k
C2 Net-_C2-Pad1_ Net-_C1-Pad1_ 1n
R2 +15V Net-_C2-Pad1_ 22k
R4 Net-_C7-Pad1_ Net-_Q2-Pad1_ 47k
C1 Net-_C1-Pad1_ IN 10u
XRV1 Net-_Q2-Pad1_ Net-_C5-Pad1_ OUT voltage_divider
R6 Net-_C2-Pad1_ Net-_C1-Pad1_ 2.2Meg
C6 Net-_C6-Pad1_ Net-_C2-Pad1_ 47n
R7 Net-_Q2-Pad1_ Net-_C6-Pad1_ 1.2Meg
C5 Net-_C5-Pad1_ Net-_C2-Pad1_ 2.2n
R8 Net-_C7-Pad1_ +15V 100k
C7 Net-_C7-Pad1_ +15V 47n
C4 GND Net-_C4-Pad2_ 10u
R5 Net-_C4-Pad2_ GND 1.5k
C3 GND Net-_C3-Pad2_ 10u
R3 Net-_C3-Pad2_ GND 1k
.end
