.title KiCad schematic
Q1 OUT_A Net-_Q1-Pad2_ Net-_Q1-Pad3_ BC547B
Q3 OUT_B Net-_Q3-Pad2_ Net-_Q1-Pad3_ BC547B
Q4 OUT_A Net-_Q4-Pad2_ Net-_Q4-Pad3_ BC547B
Q6 OUT_B Net-_Q6-Pad2_ Net-_Q4-Pad3_ BC547B
Q2 Net-_Q1-Pad3_ Net-_C1-Pad1_ Net-_Q2-Pad3_ BC547B
Q5 Net-_Q4-Pad3_ Net-_Q5-Pad2_ Net-_Q5-Pad3_ BC547B
R2 Net-_Q1-Pad2_ CV_IN 47
R12 CV_IN Net-_Q6-Pad2_ 47
R7 GND Net-_Q3-Pad2_ 47
R8 Net-_Q4-Pad2_ GND 47
R3 +15V OUT_B 680
R14 +15V OUT_A 680
R13 +15V OUT_B 680
R1 +15V OUT_A 680
R9 Net-_Q5-Pad3_ -15V 680
R6 Net-_Q2-Pad3_ -15V 680
C2 GND Net-_C2-Pad2_ 0.1u
R11 Net-_C2-Pad2_ -15V 3k
R10 +15V Net-_C2-Pad2_ 1k
C1 Net-_C1-Pad1_ NC_01 1u
R4 Net-_C2-Pad2_ Net-_C1-Pad1_ 57
R5 Net-_C2-Pad2_ Net-_Q5-Pad2_ 57
.end
