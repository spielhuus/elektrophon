.title KiCad schematic
.include diode_opamp.cir
.control
* Save only the output values
save v(OUT)
* 44100Hz sampling frequency
tran 22.675u 6
wrdata output v(OUT)
* you can use output.data as input for scripts
.endc
.subckt voltage_divider n1 n2 n3
R1 n1 n2 90kOhm
R2 n2 n3 10kOhm
.ends voltage_divider
V1 +15V 0 DC 15
V2 -15V 0 DC -15
a1 %v([IN]) filesrc

.model filesrc filesource (file="input.spice" amploffset=[0] amplscale=[5]
+                          timeoffset=0 timescale=1
+                          timerelative=false amplstep=false)

.end
