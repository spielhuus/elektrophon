.title KiCad schematic
R3 Net-_R3-Pad1_ /TRIGGER 27k
XU1 Net-_D1-Pad2_ Net-_R7-Pad2_ Net-_R3-Pad1_ +15V Net-_D2-Pad1_ Net-_D3-Pad1_ Net-_D6-Pad2_ Net-_R11-Pad1_ Net-_R11-Pad1_ Net-_C5-Pad1_ -15V Net-_R10-Pad2_ Net-_R11-Pad1_ Net-_D5-Pad1_ TL074c
R4 GND /TRIGGER 470k
R8 Net-_D1-Pad2_ Net-_R3-Pad1_ 470k
R7 GND Net-_R7-Pad2_ 27k
D2 Net-_D1-Pad1_ Net-_D2-Pad1_ D1N4148
D1 Net-_D1-Pad2_ Net-_D1-Pad1_ D1N4148
R9 Net-_R10-Pad2_ Net-_D2-Pad1_ 2.2k
R10 GND Net-_R10-Pad2_ 47k
D5 Net-_D5-Pad2_ Net-_D5-Pad1_ D1N4148
R5 Net-_D5-Pad2_ Net-_R3-Pad1_ 390k
R6 GND Net-_D5-Pad2_ 47k
D4 Net-_D3-Pad1_ Net-_D4-Pad1_ D1N4148
D3 Net-_D3-Pad2_ Net-_D3-Pad1_ D1N4148
D6 Net-_D6-Pad2_ Net-_D3-Pad2_ D1N4148
D7 Net-_D4-Pad1_ Net-_D6-Pad2_ D1N4148
C5 Net-_C5-Pad1_ GND 2.2u
D9 Net-_D9-Pad2_ Net-_D6-Pad2_ D1N4148
R11 Net-_R11-Pad1_ Net-_D3-Pad1_ 10k
D8 Net-_D6-Pad2_ Net-_D8-Pad1_ D1N4148
XRV2 Net-_C5-Pad1_ Net-_D9-Pad2_ Net-_D9-Pad2_ POT2
XRV1 Net-_C5-Pad1_ Net-_D8-Pad1_ Net-_D8-Pad1_ POT1
R12 /OUT Net-_R11-Pad1_ 2,2k
R13 GND /OUT 2.2k
.end
