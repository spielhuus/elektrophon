.title KiCad schematic
R6 Net-_R4-Pad2_ GND 36k
R4 Net-_R3-Pad2_ Net-_R4-Pad2_ 47k
R3 Net-_R2-Pad2_ Net-_R3-Pad2_ 47k
R2 Net-_R1-Pad2_ Net-_R2-Pad2_ 47k
R1 +15V Net-_R1-Pad2_ 300k
R7 Net-_R12-Pad2_ CV 47k
R8 Net-_R13-Pad2_ CV 47k
R9 Net-_R14-Pad2_ CV 47k
R10 Net-_R10-Pad1_ CV 47k
R13 Net-_Q4-Pad2_ Net-_R13-Pad2_ 750k
R14 Net-_Q2-Pad2_ Net-_R14-Pad2_ 750k
R15 Net-_Q3-Pad2_ Net-_R10-Pad1_ 750k
R12 Net-_Q1-Pad2_ Net-_R12-Pad2_ 750k
XU5 Net-_Q4-Pad3_ NC_01 INPUT_B GND Net-_R26-Pad2_ -15V NC_02 NC_03 NC_04 NC_05 +15V Net-_R25-Pad2_ GND INPUT_A NC_06 Net-_Q1-Pad3_ LM13700d
XU6 Net-_Q3-Pad3_ NC_07 INPUT_D GND Net-_R28-Pad2_ -15V NC_08 NC_09 NC_10 NC_11 +15V Net-_R27-Pad2_ GND INPUT_C NC_12 Net-_Q2-Pad3_ LM13700d
Q4 Net-_Q4-Pad1_ Net-_Q4-Pad2_ Net-_Q4-Pad3_ BC556B
D1 Net-_D1-Pad1_ +15V D1N4148
R5 Net-_D1-Pad1_ Net-_Q1-Pad1_ 33k
Q3 Net-_Q3-Pad1_ Net-_Q3-Pad2_ Net-_Q3-Pad3_ BC556B
Q2 Net-_Q2-Pad1_ Net-_Q2-Pad2_ Net-_Q2-Pad3_ BC556B
R27 NC_13 Net-_R27-Pad2_ 100k
R26 NC_14 Net-_R26-Pad2_ 100k
R25 NC_15 Net-_R25-Pad2_ 100k
R28 NC_16 Net-_R28-Pad2_ 100k
R19 Net-_Q2-Pad2_ Net-_Q3-Pad1_ 33k
R18 Net-_Q4-Pad2_ Net-_Q2-Pad1_ 33k
R17 Net-_Q1-Pad2_ Net-_Q4-Pad1_ 33k
XU1 Net-_R1-Pad2_ Net-_R12-Pad2_ +15V GND Net-_Q1-Pad2_ LT1014x_30V
XU2 Net-_R2-Pad2_ Net-_R13-Pad2_ +15V GND Net-_Q4-Pad2_ LT1014x_30V
XU3 Net-_R3-Pad2_ Net-_R14-Pad2_ +15V GND Net-_Q2-Pad2_ LT1014x_30V
XU4 Net-_R4-Pad2_ Net-_R10-Pad1_ +15V GND Net-_Q3-Pad2_ LT1014x_30V
Q1 Net-_Q1-Pad1_ Net-_Q1-Pad2_ Net-_Q1-Pad3_ BC556B
.end
