.title KiCad schematic
R1 Net-_C1-Pad2_ Net-_C2-Pad1_ 100k
XU2 GND Net-_C1-Pad2_ VP VM Net-_C1-Pad1_ TL072
R2 Net-_C1-Pad1_ Net-_C1-Pad2_ 100k
C1 Net-_C1-Pad1_ Net-_C1-Pad2_ 47p
R3 INTEGRTOR Net-_C1-Pad1_ 200k
R4 GND INTEGRTOR 10k
V1 VP GND 15
V2 VM GND -15
V3 IN_SIGNAL GND sin(0 5 1k 0 0)
Q1 Net-_Q1-Pad1_ INTEGRTOR Net-_Q1-Pad3_ BC547
Q2 Net-_Q2-Pad1_ GND Net-_Q1-Pad3_ BC547
R5 Net-_Q1-Pad1_ VP 15k
R7 Net-_Q2-Pad1_ VP 15k
R9 Net-_Q2-Pad1_ Net-_R12-Pad1_ 10k
R10 Net-_Q1-Pad1_ Net-_R10-Pad2_ 10k
R11 Net-_R10-Pad2_ GND 220k
R12 Net-_R12-Pad1_ OUT 220k
C2 Net-_C2-Pad1_ IN_SIGNAL 100n
IRV1 VP Net-_R13-Pad2_ GND dc 0 ac 0
XU4 GND Net-_R13-Pad1_ VP VM Net-_R14-Pad1_ TL072
R8 Net-_R13-Pad1_ IN_CV 68k
R13 Net-_R13-Pad1_ Net-_R13-Pad2_ 100k
R14 Net-_R14-Pad1_ Net-_R13-Pad1_ 100k
R15 Net-_Q3-Pad2_ Net-_R14-Pad1_ 22k
Q3 NC_01 Net-_Q3-Pad2_ GND BC547
R17 VM Net-_Q1-Pad3_ 15k
V4 IN_CV GND pulse(0 5 0 10m 10m 1m)
V5 NC_02 GND dc 12
R16 Net-_R16-Pad1_ Net-_Q3-Pad2_ 22k
.tran 1u 10m 
.end
