.title KiCad schematic
R11 Net-_C4-Pad1_ Net-_R11-Pad2_ 100k
R2 Net-_R11-Pad2_ Net-_R2-Pad2_ 820k
XRV5 +5V Net-_R15-Pad1_ -5V TRIM
R17 GND Net-_Q1-Pad1_ 22k
Q2 Net-_Q2-Pad3_ Net-_Q1-Pad2_ Net-_Q1-Pad1_ BC556B
Q1 Net-_Q1-Pad1_ Net-_Q1-Pad1_ Net-_Q1-Pad2_ BC556B
R14 Net-_Q1-Pad1_ Net-_R14-Pad2_ 51k
R4 Net-_R14-Pad2_ Net-_R4-Pad2_ 100k
XU2 Net-_Q1-Pad2_ Net-_R14-Pad2_ GND -15V GND Net-_C4-Pad1_ /IN +15V TL072c
R15 Net-_R15-Pad1_ Net-_R12-Pad2_ 3M
R63 /IN Net-_C4-Pad1_ 100k
C4 Net-_C4-Pad1_ /IN 47p
R12 GND Net-_R12-Pad2_ 10k
R9 GND Net-_R12-Pad2_ 100k
R3 GND Net-_R1-Pad1_ 10k
R1 Net-_R1-Pad1_ Net-_J2-PadT_ 100k
XJ2 GND Net-_J2-PadT_ NC_01 IN
R16 Net-_R16-Pad1_ Net-_Q2-Pad3_ 10k
XRV1 +5V Net-_R2-Pad2_ -5V POT
XRV2 +5V Net-_R4-Pad2_ GND POT
R6 Net-_R6-Pad1_ +5V 51k
R13 Net-_C3-Pad2_ +5V 100k
C3 -15V Net-_C3-Pad2_ 10u
R10 Net-_C4-Pad1_ Net-_R10-Pad2_ 100k
XJ3 GND Net-_J3-PadT_ NC_02 LEVEL
XRV3 Net-_J3-PadT_ Net-_R10-Pad2_ GND POT
XRV4 Net-_J1-PadT_ Net-_R5-Pad2_ GND POT
XJ1 GND Net-_J1-PadT_ NC_03 CV
R5 Net-_R14-Pad2_ Net-_R5-Pad2_ 100k
XU1 Net-_R16-Pad1_ Net-_U1-Pad12_ Net-_R1-Pad1_ Net-_R12-Pad2_ Net-_C4-Pad1_ -15V NC_04 NC_05 NC_06 NC_07 +15V Net-_U1-Pad12_ GND Net-_R6-Pad1_ Net-_R6-Pad1_ Net-_C3-Pad2_ LM13700d
.end
