.title KiCad schematic
XU1 IN_Xa IN_Xa GND -15V GND IN_Ya IN_Ya +15V TL072c
XU2 OUT_a Net-_R1-Pad1_ Net-_U2-Pad3_ -15V GND IN_Za IN_Za +15V TL072c
XU3 IN_Xa GND IN_Ya GND -15V IN_Za Net-_U2-Pad3_ +15V AD633
R2 OUT_a Net-_R1-Pad1_ 10k
R1 Net-_R1-Pad1_ GND 10k
.end
