.title KiCad schematic
C11 Net-_C11-Pad1_ GND 22n
C12 Net-_C1-Pad1_ Net-_C12-Pad2_ 220n
R24 Net-_C12-Pad2_ NC_01 15k
R25 Net-_C11-Pad1_ Net-_C12-Pad2_ 15k
Q1 Net-_Q1-Pad1_ Net-_Q1-Pad2_ Net-_C1-Pad1_ BC846B
Q2 Net-_C1-Pad1_ Net-_Q1-Pad1_ +15V BC556B
R1 Net-_Q1-Pad2_ Net-_C11-Pad1_ 10k
R2 GND Net-_C1-Pad1_ 1.5k
R3 /OUT GND 10k
C1 Net-_C1-Pad1_ /OUT 100u
.end
