.title KiCad schematic
XU1 Net-_C1-Pad1_ Net-_C3-Pad2_ +15V GND 4069UB
R2 Net-_C2-Pad2_ Net-_C1-Pad1_ 100k
R1 Net-_C1-Pad2_ NC_01 100k
C3 /OUT Net-_C3-Pad2_ 10u
R6 GND /OUT 1k
C1 Net-_C1-Pad1_ Net-_C1-Pad2_ 22n
R3 Net-_C3-Pad2_ Net-_C2-Pad2_ 100k
C2 GND Net-_C2-Pad2_ 1.8n
.end
