.title KiCad schematic
.include ../../../lib/spice/opamp/TL072.lib
.include ../../../lib/spice/diode/1N4148.mod
.include 'Overdrive 250.cir'
.control
* Save only the output values
save v(OUT)
* 44100Hz sampling frequency
tran 22.675u 6
wrdata build/output v(OUT)
* you can use output.data as input for scripts
.endc
.subckt voltage_divider n1 n2 n3
R1 n1 n2 499kOhm
R2 n2 n3 1kOhm
.ends voltage_divider

V1 +5V 0 DC 5
a1 %v([IN]) filesrc

.model filesrc filesource (file="build/input.spice" amploffset=[0] amplscale=[5]
+                          timeoffset=0 timescale=1
+                          timerelative=false amplstep=false)

.end
.measure tran ymax MAX v(OUT) from=0m to=30m
.measure tran ymax RMS v(OUT) from=0m to=30m

