.title KiCad schematic
XU1 Net-_R2-Pad1_ Net-_C3-Pad1_ +15V GND Net-_C4-Pad1_ TL072
R4 +15V Net-_C2-Pad1_ 22k
R5 Net-_C2-Pad1_ GND 220k
R1 Net-_C1-Pad2_ GND 25k
R2 Net-_R2-Pad1_ Net-_C1-Pad1_ 10k
R6 Net-_C2-Pad1_ Net-_R2-Pad1_ 470k
C1 Net-_C1-Pad1_ Net-_C1-Pad2_ 10n
C2 Net-_C2-Pad1_ GND 10u
C4 Net-_C4-Pad1_ Net-_C3-Pad1_ 22p
R7 Net-_C4-Pad1_ Net-_C3-Pad1_ 1Meg
C3 Net-_C3-Pad1_ Net-_C3-Pad2_ 4.7n
R3 Net-_C3-Pad2_ Net-_R3-Pad2_ 4.7k
XRV1 GND GND Net-_R3-Pad2_ voltage_divider
C5 Net-_C4-Pad1_ Net-_C5-Pad2_ 4.7u
R8 OUT Net-_C5-Pad2_ 10k
D1 GND OUT D1N4148
D2 OUT Net-_D2-Pad2_ D1N4148
D3 Net-_D2-Pad2_ GND D1N4148
C6 GND OUT 1n
R9 IN Net-_C1-Pad2_ 100k
.end
