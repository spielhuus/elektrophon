.title KiCad schematic
V1 +15V GND +15
V2 -15V GND -15
Q1 OUT_A Net-_C5-Pad1_ Net-_Q1-Pad3_ BC547B
Q3 OUT_B Net-_Q3-Pad2_ Net-_Q1-Pad3_ BC547B
Q4 OUT_A Net-_Q3-Pad2_ Net-_Q4-Pad3_ BC547B
Q6 OUT_B Net-_C5-Pad1_ Net-_Q4-Pad3_ BC547B
R9 +15V OUT_A 270
R13 +15V OUT_B 270
Q2 Net-_Q1-Pad3_ Net-_C6-Pad1_ Net-_Q2-Pad3_ BC547B
Q5 Net-_Q4-Pad3_ Net-_Q5-Pad2_ Net-_Q2-Pad3_ BC547B
R16 +15V Net-_C7-Pad2_ 4.7k
R17 Net-_C7-Pad2_ Net-_C9-Pad1_ 3.3k
R18 Net-_C9-Pad1_ GND 2.2k
C8 Net-_C7-Pad2_ GND 0.1u
C9 Net-_C9-Pad1_ GND 0.1u
V3 +5V GND dc 5
R15 Net-_C7-Pad2_ Net-_C5-Pad1_ 2.2k
R11 Net-_C7-Pad2_ Net-_Q3-Pad2_ 2.2k
R14 Net-_C9-Pad1_ Net-_Q5-Pad2_ 2.2k
R10 Net-_C9-Pad1_ Net-_C6-Pad1_ 2.2k
C7 GND Net-_C7-Pad2_ 0.1u
C5 Net-_C5-Pad1_ in 0.1u
C6 Net-_C6-Pad1_ cv 0.1u
R12 Net-_Q2-Pad3_ GND 270
XU1 Net-_R3-Pad1_ Net-_R1-Pad1_ GND -15V GND Net-_R2-Pad1_ Net-_R4-Pad1_ +15V OPA2134d
R3 Net-_R3-Pad1_ Net-_R1-Pad1_ 100k
R5 Net-_R5-Pad1_ Net-_R3-Pad1_ 100k
R1 Net-_R1-Pad1_ Net-_R1-Pad2_ 100k
XRV1 GND Net-_R1-Pad2_ Net-_J1-PadT_ voltage_divider_1
VJ1 Net-_J1-PadT_ GND dc 5 sin(0 20m 1k)
VJ2 Net-_J2-PadT_ GND dc 5 sin(0 20m 200)
XRV2 GND Net-_R2-Pad2_ Net-_J2-PadT_ voltage_divider_1
R2 Net-_R2-Pad1_ Net-_R2-Pad2_ 100k
R4 Net-_R4-Pad1_ Net-_R2-Pad1_ 100k
R6 Net-_R6-Pad1_ Net-_R4-Pad1_ 100k
R8 GND Net-_R6-Pad1_ 1k
R7 GND Net-_R5-Pad1_ 1k
XU2 Net-_R19-Pad1_ Net-_R19-Pad1_ Net-_R5-Pad1_ -15V Net-_R6-Pad1_ Net-_R20-Pad1_ Net-_R20-Pad1_ +15V OPA2134d
R19 Net-_R19-Pad1_ in 2.2k
R20 Net-_R20-Pad1_ cv 2.2k
.end
