.title KiCad schematic
XU1 Net-_C1-Pad2_ Net-_C1-Pad1_ +5V GND 4069UB
R2 Net-_C1-Pad1_ Net-_C1-Pad2_ 100k
R1 Net-_C1-Pad2_ IN 100k
C1 Net-_C1-Pad1_ Net-_C1-Pad2_ 0.01u
C3 OUT Net-_C1-Pad1_ 1u
R3 GND OUT 100k
.end
