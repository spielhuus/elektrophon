.title KiCad schematic
XRV2 CV_B Net-_R16-Pad2_ CV_A voltage_divider_2
R16 CV_IN Net-_R16-Pad2_ 100k
XU1 Net-_C1-Pad1_ CV_B GND -15V GND CV_A CV +15V TL072c
R12 CV_B OFFSET 200k
R14 CV_A Net-_C1-Pad1_ 100k
C2 CV CV_A 100n
C1 Net-_C1-Pad1_ CV_B 100n
R15 CV CV_A 33k
R13 Net-_C1-Pad1_ CV_B 100k
R1 Net-_Q2-Pad2_ GND 6.8k
Q1 Net-_Q1-Pad2_ Net-_Q1-Pad2_ +15V q2n3906
Q2 Net-_Q2-Pad2_ Net-_Q2-Pad2_ Net-_Q1-Pad2_ q2n3906
R11 +15V Net-_Q8-Pad1_ 1k
R2 +15V Net-_R2-Pad2_ 100
XRV1 Net-_R2-Pad2_ Net-_Q3-Pad1_ Net-_Q3-Pad1_ voltage_divider_1
D6 Net-_D6-Pad2_ Net-_D6-Pad1_ D1N4148
R9 Net-_D6-Pad2_ Net-_D4-Pad2_ 100
R6 Net-_D4-Pad2_ CV 100
R7 GND Net-_D3-Pad2_ 100
R4 Net-_D3-Pad2_ Net-_D1-Pad2_ 100
D4 Net-_D4-Pad2_ Net-_D4-Pad1_ D1N4148
D2 CV Net-_D2-Pad1_ D1N4148
D5 GND Net-_D4-Pad1_ D1N4148
D3 Net-_D3-Pad2_ Net-_D2-Pad1_ D1N4148
R10 Net-_D6-Pad1_ -15V 1meg
R8 Net-_D4-Pad1_ -15V 1meg
R5 Net-_D2-Pad1_ -15V 1meg
D1 Net-_D1-Pad2_ Net-_D1-Pad1_ D1N4148
R3 Net-_D1-Pad1_ -15V 1meg
Q4 I1 Net-_D1-Pad1_ Net-_Q4-Pad1_ q2n3906
Q5 I2 Net-_D2-Pad1_ Net-_Q4-Pad1_ q2n3906
Q6 I3 Net-_D4-Pad1_ Net-_Q4-Pad1_ q2n3906
Q9 I4 Net-_D6-Pad1_ Net-_Q4-Pad1_ q2n3906
Q8 Net-_Q4-Pad1_ Net-_Q2-Pad2_ Net-_Q8-Pad1_ q2n3906
Q7 Net-_D6-Pad2_ Net-_Q2-Pad2_ Net-_Q3-Pad1_ q2n3906
Q3 Net-_D1-Pad2_ Net-_Q2-Pad2_ Net-_Q3-Pad1_ q2n3906
.end
