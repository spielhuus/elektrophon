.title KiCad schematic
XU3 Net-_C5-Pad2_ Net-_C6-Pad1_ +15V -15V Net-_C6-Pad1_ TL072
C6 Net-_C6-Pad1_ Net-_C6-Pad2_ 47n
R6 Net-_C5-Pad2_ Net-_C6-Pad2_ 15k
R5 Net-_C6-Pad2_ NC_01 15k
C5 GND Net-_C5-Pad2_ 4.7n
XU4 Net-_C8-Pad1_ /OUT +15V -15V /OUT TL072
C7 Net-_C7-Pad1_ Net-_C6-Pad1_ 47n
R8 /OUT Net-_C7-Pad1_ 4.7k
R7 GND Net-_C8-Pad1_ 40k
C8 Net-_C8-Pad1_ Net-_C7-Pad1_ 47n
.end
