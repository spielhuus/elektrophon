.title KiCad schematic
XU1 OUT Net-_C2-Pad1_ +5V GND CD4069UB
R3 OUT Net-_C2-Pad1_ 1Meg
XU2 Net-_R2-Pad1_ Net-_R1-Pad1_ GND -15V NC_01 NC_02 NC_03 +15V TL072c
C1 Net-_C1-Pad1_ IN 0.22u
R1 Net-_R1-Pad1_ Net-_C1-Pad1_ 100k
R2 Net-_R2-Pad1_ Net-_R1-Pad1_ 100k
R4 Net-_C2-Pad2_ Net-_R2-Pad1_ 10k
C2 Net-_C2-Pad1_ Net-_C2-Pad2_ 22n
.end
