.title KiCad schematic
XU1 Net-_R12-Pad1_ Net-_R1-Pad1_ +15V -15V Net-_D2-Pad2_ TL072
R1 Net-_R1-Pad1_ CV_IN 100k
R13 Net-_D2-Pad2_ Net-_R1-Pad1_ 62k
Q7 Net-_D6-Pad2_ Net-_Q2-Pad2_ Net-_Q3-Pad1_ q2n3906
Q8 Net-_Q4-Pad1_ Net-_Q2-Pad2_ Net-_Q8-Pad1_ q2n3906
Q9 Net-_Q9-Pad3_ Net-_D6-Pad1_ Net-_Q4-Pad1_ q2n3906
Q6 Net-_Q6-Pad3_ Net-_D4-Pad1_ Net-_Q4-Pad1_ q2n3906
Q5 Net-_Q5-Pad3_ Net-_D2-Pad1_ Net-_Q4-Pad1_ q2n3906
Q4 Net-_Q4-Pad3_ Net-_D1-Pad1_ Net-_Q4-Pad1_ q2n3906
R3 Net-_D1-Pad1_ -15V 1meg
D1 Net-_D1-Pad2_ Net-_D1-Pad1_ D1N4148
R5 Net-_D2-Pad1_ -15V 1meg
R8 Net-_D4-Pad1_ -15V 1meg
R10 Net-_D6-Pad1_ -15V 1meg
D3 Net-_D3-Pad2_ Net-_D2-Pad1_ D1N4148
D5 GND Net-_D4-Pad1_ D1N4148
D2 Net-_D2-Pad2_ Net-_D2-Pad1_ D1N4148
D4 Net-_D4-Pad2_ Net-_D4-Pad1_ D1N4148
R4 Net-_D3-Pad2_ Net-_D1-Pad2_ 100
R7 GND Net-_D3-Pad2_ 100
R6 Net-_D4-Pad2_ Net-_D2-Pad2_ 100
R9 Net-_D6-Pad2_ Net-_D4-Pad2_ 100
D6 Net-_D6-Pad2_ Net-_D6-Pad1_ D1N4148
XRV1 Net-_R2-Pad2_ Net-_Q3-Pad1_ Net-_Q3-Pad1_ voltage_divider_1
R2 +15V Net-_R2-Pad2_ 100
R11 +15V Net-_Q8-Pad1_ 1k
R12 Net-_R12-Pad1_ GND 39k
R16 Net-_Q4-Pad3_ GND 220
R17 Net-_Q5-Pad3_ GND 220
R18 Net-_Q6-Pad3_ GND 220
R19 Net-_Q9-Pad3_ GND 220
Q1 Net-_Q1-Pad2_ Net-_Q1-Pad2_ +15V q2n3906
Q2 Net-_Q2-Pad2_ Net-_Q2-Pad2_ Net-_Q1-Pad2_ q2n3906
R14 Net-_Q2-Pad2_ GND 6.8k
Q3 Net-_D1-Pad2_ Net-_Q2-Pad2_ Net-_Q3-Pad1_ q2n3906
.end
