.title KiCad schematic
XU1 Net-_R1-Pad1_ Net-_R2-Pad1_ +5V GND 4069UB
R2 Net-_R2-Pad1_ Net-_R1-Pad1_ 10k
R3 Net-_C1-Pad2_ Net-_R2-Pad1_ 20k
XU2 Net-_C1-Pad2_ Net-_C1-Pad1_ +5V GND 4069UB
XU3 Net-_C2-Pad2_ OUT +5V GND 4069UB
C2 OUT Net-_C2-Pad2_ 0.01u
XRV1 NC_01 Net-_R4-Pad1_ OUT voltage_divider_1
R1 Net-_R1-Pad1_ IN 10k
C1 Net-_C1-Pad1_ Net-_C1-Pad2_ 0.1u
R5 Net-_C2-Pad2_ Net-_C1-Pad1_ 20k
R4 Net-_R4-Pad1_ Net-_C1-Pad2_ 6.8k
.end
