.title KiCad schematic
R4 Net-_C7-Pad2_ Net-_C3-Pad1_ 1Meg
XRV1 Net-_R3-Pad1_ Net-_RV1-Pad2_ Net-_R7-Pad2_ voltage_divider_1
R3 Net-_R3-Pad1_ Net-_R2-Pad2_ 100k
R1 GND Net-_C2-Pad2_ 10k
R2 Net-_C1-Pad1_ Net-_R2-Pad2_ 100k
C1 Net-_C1-Pad1_ Net-_C1-Pad2_ 100n
C3 Net-_C3-Pad1_ Net-_C3-Pad2_ 470n
XU1 Net-_R5-Pad2_ Net-_C1-Pad2_ Net-_R2-Pad2_ Net-_RV1-Pad2_ Net-_C3-Pad1_ Net-_C7-Pad2_ GND NC_01 +5V Net-_C8-Pad1_ Net-_R11-Pad1_ NC_02 +5V +5V CD4069UBhex
C2 Net-_C2-Pad1_ Net-_C2-Pad2_ 10n
R5 Net-_C2-Pad1_ Net-_R5-Pad2_ 470k
R6 Net-_R5-Pad2_ Net-_C1-Pad2_ 470k
R7 Net-_C3-Pad2_ Net-_R7-Pad2_ 10k
D2 Net-_C3-Pad1_ Net-_D2-Pad2_ D1N4148
D1 Net-_D1-Pad1_ Net-_C3-Pad1_ D1N4148
C7 Net-_C7-Pad1_ Net-_C7-Pad2_ 100n
R11 Net-_R11-Pad1_ Net-_C7-Pad1_ 100k
R13 Net-_C8-Pad1_ Net-_R11-Pad1_ 1Meg
C8 Net-_C8-Pad1_ OUT 10u
R14 GND OUT 10k
R8 Net-_R11-Pad1_ Net-_C1-Pad2_ 100k
D6 Net-_D4-Pad2_ Net-_C7-Pad2_ D1N4148
D4 Net-_D2-Pad2_ Net-_D4-Pad2_ D1N4148
D5 Net-_C7-Pad2_ Net-_D3-Pad1_ D1N4148
D3 Net-_D3-Pad1_ Net-_D1-Pad1_ D1N4148
R9 IN Net-_C2-Pad2_ 100k
.end
