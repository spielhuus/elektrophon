.title KiCad schematic
XU1 Net-_R2-Pad2_ SAW_IN GND -15V Net-_R1-Pad1_ Net-_R3-Pad2_ OUT +15V TL072c
R1 Net-_R1-Pad1_ SAW_IN 49.9k
R2 Net-_R1-Pad1_ Net-_R2-Pad2_ 300k
R4 OUT Net-_R3-Pad2_ 100k
R3 GND Net-_R3-Pad2_ 49.9k
.end
