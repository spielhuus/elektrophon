.title KiCad schematic
R58 Net-_C1-Pad1_ Net-_R57-Pad1_ 100k
C1 Net-_C1-Pad1_ GND 22u
XU6 +5V Net-_C2-Pad2_ Net-_C1-Pad1_ -15V GND Net-_C3-Pad2_ -5V +15V TL072c
R61 Net-_C3-Pad2_ +5V 100k
R57 Net-_R57-Pad1_ +15V 10k
R60 +5V Net-_C2-Pad2_ 100k
C2 +5V Net-_C2-Pad2_ 22u
R59 GND Net-_C2-Pad2_ 100k
R62 -5V Net-_C3-Pad2_ 100k
C3 -5V Net-_C3-Pad2_ 22u
XU7 Net-_R57-Pad1_ GND Net-_R57-Pad1_ TL431
.end
