.title KiCad schematic
XU2 Net-_C9-Pad2_ Net-_R15-Pad1_ Net-_R16-Pad1_ -15V GND Net-_U2-Pad6_ Net-_U2-Pad6_ +15V TL072c
R14 /IN GND 100k
R18 GND Net-_R16-Pad1_ 2.7k
R16 Net-_R16-Pad1_ +15V 22k
R15 Net-_R15-Pad1_ /IN 10k
R17 Net-_C9-Pad2_ Net-_R16-Pad1_ 1Meg
C9 Net-_C9-Pad1_ Net-_C9-Pad2_ 560p
R19 +15V Net-_C9-Pad1_ 56k
C10 Net-_C10-Pad1_ GND 0.01u
XU3 GND Net-_C9-Pad1_ Net-_C11-Pad2_ +15V Net-_C10-Pad1_ Net-_C12-Pad1_ Net-_C12-Pad1_ +15V TLC555
XU4 GND Net-_C11-Pad1_ Net-_R22-Pad2_ Net-_C11-Pad1_ Net-_C13-Pad1_ Net-_C14-Pad1_ Net-_C14-Pad1_ +15V TLC555
XRV3 Net-_R20-Pad1_ Net-_R20-Pad1_ +15V POT1
R20 Net-_R20-Pad1_ Net-_C12-Pad1_ 1k
C12 Net-_C12-Pad1_ GND 2.2u
C11 Net-_C11-Pad1_ Net-_C11-Pad2_ 560p
R21 +15V Net-_C11-Pad1_ 56k
C13 Net-_C13-Pad1_ GND 0.01u
XRV4 Net-_R23-Pad1_ Net-_R23-Pad1_ +15V POT2
R23 Net-_R23-Pad1_ Net-_C14-Pad1_ 1k
C14 Net-_C14-Pad1_ GND 2.2u
R22 /del_out Net-_R22-Pad2_ 2.7k
R24 GND /del_out 1.8k
.end
