.title KiCad schematic
Q1 OUT_A CV_IN Net-_Q1-Pad3_ BC547B
Q3 OUT_B GND Net-_Q1-Pad3_ BC547B
Q4 OUT_A GND Net-_Q4-Pad3_ BC547B
Q6 OUT_B CV_IN Net-_Q4-Pad3_ BC547B
Q2 Net-_Q1-Pad3_ Net-_C1-Pad1_ Net-_Q2-Pad3_ BC547B
Q5 Net-_Q4-Pad3_ Net-_Q5-Pad2_ Net-_Q2-Pad3_ BC547B
R3 +15V OUT_B 720
R1 +15V OUT_A 720
R7 Net-_R2-Pad2_ OUT 440k
R6 GND Net-_R5-Pad2_ 440k
XU1 Net-_R5-Pad2_ Net-_R2-Pad2_ +15V -15V OUT TL072
R2 OUT_A Net-_R2-Pad2_ 10k
R5 OUT_B Net-_R5-Pad2_ 10k
R8 Net-_Q2-Pad3_ -15V 720
C1 Net-_C1-Pad1_ AUDIO_IN 0.22u
R11 Net-_C2-Pad2_ -15V 1k
R10 +15V Net-_C2-Pad2_ 3k
R9 Net-_C2-Pad2_ Net-_Q5-Pad2_ 2.2k
R4 Net-_C2-Pad2_ Net-_C1-Pad1_ 2.2k
C2 GND Net-_C2-Pad2_ 0.1u
.end
