.title KiCad schematic
XU5 Net-_C9-Pad2_ Net-_C10-Pad1_ +15V -15V Net-_C10-Pad1_ TL072
C10 Net-_C10-Pad1_ Net-_C10-Pad2_ 10n
R10 Net-_C9-Pad2_ Net-_C10-Pad2_ 15k
R9 Net-_C10-Pad2_ NC_01 15k
C9 GND Net-_C9-Pad2_ 910p
XU6 Net-_C12-Pad1_ /OUT +15V -15V /OUT TL072
C11 Net-_C11-Pad1_ Net-_C10-Pad1_ 10n
R12 /OUT Net-_C11-Pad1_ 4.7k
R11 GND Net-_C12-Pad1_ 40k
C12 Net-_C12-Pad1_ Net-_C11-Pad1_ 10n
.end
