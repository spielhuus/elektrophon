.title KiCad schematic
XU1 Net-_C4-Pad1_ Net-_C2-Pad1_ +15V GND 4069UB
C1 Net-_C1-Pad1_ Net-_C1-Pad2_ 22n
C3 /OUT Net-_C2-Pad1_ 10u
R6 GND /OUT 1k
C2 Net-_C2-Pad1_ Net-_C1-Pad1_ 22n
R3 GND Net-_C1-Pad1_ 10
R1 Net-_C5-Pad2_ Net-_C4-Pad1_ 100k
R4 Net-_C2-Pad1_ Net-_C5-Pad2_ 100k
C5 GND Net-_C5-Pad2_ 22n
C4 Net-_C4-Pad1_ Net-_C1-Pad2_ 100n
R2 Net-_C1-Pad2_ NC_01 10k
.end
