.title KiCad schematic
XU1 Net-_R2-Pad1_ Net-_C2-Pad2_ Net-_R4-Pad1_ Net-_RV1-Pad2_ Net-_C3-Pad1_ Net-_C4-Pad2_ GND Net-_C6-Pad1_ Net-_C6-Pad2_ Net-_C9-Pad2_ Net-_R11-Pad1_ GND GND +5V CD4069UBhex
R1 IN GND 1Meg
R2 Net-_R2-Pad1_ Net-_C1-Pad1_ 470k
R3 Net-_C2-Pad2_ Net-_R2-Pad1_ 470k
R4 Net-_R4-Pad1_ Net-_C2-Pad1_ 100k
C1 Net-_C1-Pad1_ IN 10n
C2 Net-_C2-Pad1_ Net-_C2-Pad2_ 2.2n
R5 Net-_R5-Pad1_ Net-_R4-Pad1_ 100k
XRV1 Net-_R5-Pad1_ Net-_RV1-Pad2_ Net-_R6-Pad2_ voltage_divider_1
R6 Net-_C3-Pad2_ Net-_R6-Pad2_ 10k
C3 Net-_C3-Pad1_ Net-_C3-Pad2_ 470n
R7 Net-_C4-Pad2_ Net-_C3-Pad1_ 1Meg
D2 Net-_C3-Pad1_ Net-_C4-Pad2_ D1N4148
D1 Net-_C4-Pad2_ Net-_C3-Pad1_ D1N4148
R8 Net-_C5-Pad2_ Net-_C4-Pad1_ 100k
C4 Net-_C4-Pad1_ Net-_C4-Pad2_ 100n
C5 GND Net-_C5-Pad2_ 1.5n
R9 Net-_R9-Pad1_ Net-_C5-Pad2_ 10k
XRV2 Net-_C6-Pad2_ Net-_C6-Pad2_ Net-_R9-Pad1_ voltage_divider_2
C6 Net-_C6-Pad1_ Net-_C6-Pad2_ 150p
R10 Net-_C6-Pad1_ Net-_C5-Pad2_ 100k
R11 Net-_R11-Pad1_ Net-_C7-Pad1_ 100k
C7 Net-_C7-Pad1_ Net-_C6-Pad1_ 100n
R13 Net-_C9-Pad2_ Net-_R11-Pad1_ 220k
C9 OUT Net-_C9-Pad2_ 100n
C8 Net-_C8-Pad1_ Net-_C2-Pad2_ 100n
R12 Net-_R11-Pad1_ Net-_C8-Pad1_ 100k
R14 GND OUT 1k
.end
