.title KiCad schematic
.include "/home/etienne/Documents/elektrophon/lib/spice/opamp/TL072.lib"
.include "/home/etienne/Documents/elektrophon/lib/spice/opamp/ad633.lib"
XU1 Net-_R7-Pad1_ GND Net-_R4-Pad1_ GND -15V GND Net-_R5-Pad2_ +15V AD633
R1 NC_01 Net-_R1-Pad2_ 1k
XU2 GND Net-_R3-Pad1_ +15V -15V Net-_R7-Pad1_ TL072
R2 Net-_R2-Pad1_ Y1 100k
R4 Net-_R4-Pad1_ Net-_R2-Pad1_ 100k
XU3 GND Net-_R5-Pad1_ +15V -15V Net-_R1-Pad2_ TL072
R5 Net-_R5-Pad1_ Net-_R5-Pad2_ 100k
XU4 GND Net-_R2-Pad1_ +15V -15V Net-_R4-Pad1_ TL072
R6 Net-_R1-Pad2_ Net-_R5-Pad1_ 100k
V4 Y1 GND pulse(0 10 0 0 500m 100u 600m)
V5 NC_02 GND dc 5 sin(0 5 100)
V3 X1 GND sin(0 5 440)
V2 -15V GND -15
V1 +15V GND +15
R3 Net-_R3-Pad1_ X1 100k
R7 Net-_R7-Pad1_ Net-_R3-Pad1_ 100k
.tran 10u 20m 0 
.end
